module Adder(input wire [31:0] num0, num1, output wire [31:0] out);
    assign out = num0 + num1;
endmodule